constant PACKET : std_logic_vector(791 downto 0) :=
x"00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00" &
x"00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00" &
x"00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00" &
x"00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00" &
x"00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00" &
x"05_7e_94_9a_07_e8_81_86_c6_49_bb_eb_0a_97_40_c5_e0_19_82_ad" &
x"e7_12_f9_ec_3d_3a_57_ce_85_ad_f7_fc_3e_2b_43_d7_d8_9f_90_d3" &
x"00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00" &
x"00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00" &
x"00_00_00_00_00_00_00_00_00_00_00_00_00_00_01";
