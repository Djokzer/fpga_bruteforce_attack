��c o n s t a n t   P A C K E T   :   s t d _ l o g i c _ v e c t o r ( 8 2 3   d o w n t o   0 )   : =  
 x " 0 2 _ 6 3 _ 0 2 _ 0 5 _ 0 1 _ 0 1 _ 2 8 _ e 0 _ c 5 _ 4 0 _ 9 7 _ 0 a _ e b _ b b _ 4 9 _ c 6 _ 8 6 _ 8 1 _ e 8 _ 0 7 "   &  
 x " 9 a _ 9 4 _ 7 e _ d 3 _ 9 0 _ 9 f _ d 8 _ d 7 _ 4 3 _ 2 b _ 3 e _ f c _ f 7 _ a d _ 8 5 _ c e _ 5 7 _ 3 a _ 3 d _ e c "   &  
 x " f 9 _ 1 2 _ e 7 _ a d _ 8 2 _ 1 9 _ 0 1 _ 0 1 _ 0 1 _ 0 1 _ 0 1 _ 0 1 _ 0 1 _ 0 1 _ 0 1 _ 0 1 _ 0 1 _ 0 1 _ 0 1 _ 0 1 "   &  
 x " 0 1 _ 0 1 _ 0 1 _ 0 1 _ 0 1 _ 0 1 _ 0 1 _ 0 1 _ 0 1 _ 0 1 _ 0 1 _ 0 1 _ 0 1 _ 0 1 _ 0 1 _ 0 1 _ 0 1 _ 0 1 _ 0 1 _ 0 1 "   &  
 x " 0 1 _ 0 1 _ 0 1 _ 0 1 _ 0 1 _ 0 1 _ 0 1 _ 0 1 _ 0 1 _ 0 1 _ 0 1 _ 0 1 _ 0 1 _ 0 1 _ 0 1 _ 0 1 _ 0 1 _ 0 1 _ 0 1 _ 0 3 "   &  
 x " 0 1 _ c 0 _ 0 0 " ;  
 