library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_textio.all;
use ieee.numeric_std.all;

package pkg_sbox_init is
    constant SBOX01_INIT_VEC : std_logic_vector(16383 downto 0) :=
    x"D1310BA6_98DFB5AC_2FFD72DB_D01ADFB7_B8E1AFED_6A267E96" &
    x"BA7C9045_F12C7F99_24A19947_B3916CF7_0801F2E2_858EFC16" &
    x"636920D8_71574E69_A458FEA3_F4933D7E_0D95748F_728EB658" &
    x"718BCD58_82154AEE_7B54A41D_C25A59B5_9C30D539_2AF26013" &
    x"C5D1B023_286085F0_CA417918_B8DB38EF_8E79DCB0_603A180E" &
    x"6C9E0E8B_B01E8A3E_D71577C1_BD314B27_78AF2FDA_55605C60" &
    x"E65525F3_AA55AB94_57489862_63E81440_55CA396A_2AAB10B6" &
    x"B4CC5C34_1141E8CE_A15486AF_7C72E993_B3EE1411_636FBC2A" &
    x"2BA9C55D_741831F6_CE5C3E16_9B87931E_AFD6BA33_6C24CF5C" &
    x"7A325381_28958677_3B8F4898_6B4BB9AF_C4BFE81B_66282193" &
    x"61D809CC_FB21A991_487CAC60_5DEC8032_EF845D5D_E98575B1" &
    x"DC262302_EB651B88_23893E81_D396ACC5_0F6D6FF3_83F44239" &
    x"2E0B4482_A4842004_69C8F04A_9E1F9B5E_21C66842_F6E96C9A" &
    x"670C9C61_ABD388F0_6A51A0D2_D8542F68_960FA728_AB5133A3" &
    x"6EEF0B6C_137A3BE4_BA3BF050_7EFB2A98_A1F1651D_39AF0176" &
    x"66CA593E_82430E88_8CEE8619_456F9FB4_7D84A5C3_3B8B5EBE" &
    x"E06F75D8_85C12073_401A449F_56C16AA6_4ED3AA62_363F7706" &
    x"1BFEDF72_429B023D_37D0D724_D00A1248_DB0FEAD3_49F1C09B" &
    x"075372C9_80991B7B_25D479D8_F6E8DEF7_E3FE501A_B6794C3B" &
    x"976CE0BD_04C006BA_C1A94FB6_409F60C4_5E5C9EC2_196A2463" &
    x"68FB6FAF_3E6C53B5_1339B2EB_3B52EC6F_6DFC511F_9B30952C" &
    x"CC814544_AF5EBD09_BEE3D004_DE334AFD_660F2807_192E4BB3" &
    x"C0CBA857_45C8740F_D20B5F39_B9D3FBDB_5579C0BD_1A60320A" &
    x"D6A100C6_402C7279_679F25FE_FB1FA3CC_8EA5E9F8_DB3222F8" &
    x"3C7516DF_FD616B15_2F501EC8_AD0552AB_323DB5FA_FD238760" &
    x"53317B48_3E00DF82_9E5C57BB_CA6F8CA0_1A87562E_DF1769DB" &
    x"D542A8F6_287EFFC3_AC6732C6_8C4F5573_695B27B0_BBCA58C8" &
    x"E1FFA35D_B8F011A0_10FA3D98_FD2183B8_4AFCB56C_2DD1D35B" &
    x"9A53E479_B6F84565_D28E49BC_4BFB9790_E1DDF2DA_A4CB7E33" &
    x"62FB1341_CEE4C6E8_EF20CADA_36774C01_D07E9EFE_2BF11FB4" &
    x"95DBDA4D_AE909198_EAAD8E71_6B93D5A0_D08ED1D0_AFC725E0" &
    x"8E3C5B2F_8E7594B7_8FF6E2FB_F2122B64_8888B812_900DF01C" &
    x"4FAD5EA0_688FC31C_D1CFF191_B3A8C1AD_2F2F2218_BE0E1777" &
    x"EA752DFE_8B021FA1_E5A0CC0F_B56F74E8_18ACF3D6_CE89E299" &
    x"B4A84FE0_FD13E0B7_7CC43B81_D2ADA8D9_165FA266_80957705" &
    x"93CC7314_211A1477_E6AD2065_77B5FA86_C75442F5_FB9D35CF" &
    x"EBCDAF0C_7B3E89A0_D6411BD3_AE1E7E49_00250E2D_2071B35E" &
    x"226800BB_57B8E0AF_2464369B_F009B91E_5563911D_59DFA6AA" &
    x"78C14389_D95A537F_207D5BA2_02E5B9C5_83260376_6295CFA9" &
    x"11C81968_4E734A41_B3472DCA_7B14A94A_1B510052_9A532915" &
    x"D60F573F_BC9BC6E4_2B60A476_81E67400_08BA6FB5_571BE91F" &
    x"F296EC6B_2A0DD915_B6636521_E7B9F9B6_FF34052E_C5855664" &
    x"53B02D5D_A99F8FA1_08BA4799_6E85076A_4B7A70E9_B5B32944" &
    x"DB75092E_C4192623_AD6EA6B0_49A7DF7D_9CEE60B8_8FEDB266" &
    x"ECAA8C71_699A17FF_5664526C_C2B19EE1_193602A5_75094C29" &
    x"A0591340_E4183A3E_3F54989A_5B429D65_6B8FE4D6_99F73FD6" &
    x"A1D29C07_EFE830F5_4D2D38E6_F0255DC1_4CDD2086_8470EB26" &
    x"6382E9C6_021ECC5E_09686B3F_3EBAEFC9_3C971814_6B6A70A1" &
    x"687F3584_52A0E286_B79C5305_AA500737_3E07841C_7FDEAE5C" &
    x"8E7D44EC_5716F2B8_B03ADA37_F0500C0D_F01C1F04_0200B3FF" &
    x"AE0CF51A_3CB574B2_25837A58_DC0921BD_D19113F9_7CA92FF6" &
    x"94324773_22F54701_3AE5E581_37C2DADC_C8B57634_9AF3DDA7" &
    x"A9446146_0FD0030E_ECC8C73E_A4751E41_E238CD99_3BEA0E2F" &
    x"3280BBA1_183EB331_4E548B38_4F6DB908_6F420D03_F60A04BF" &
    x"2CB81290_24977C79_5679B072_BCAF89AF_DE9A771F_D9930810" &
    x"B38BAE12_DCCF3F2E_5512721F_2E6B7124_501ADDE6_9F84CD87" &
    x"7A584718_7408DA17_BC9F9ABC_E94B7D8C_EC7AEC3A_DB851DFA" &
    x"63094366_C464C3D2_EF1C1847_3215D908_DD433B37_24C2BA16" &
    x"12A14D43_2A65C451_50940002_133AE4DD_71DFF89E_10314E55" &
    x"81AC77D6_5F11199B_043556F1_D7A3C76B_3C11183B_5924A509" &
    x"F28FE6ED_97F1FBFA_9EBABF2C_1E153C6E_86E34570_EAE96FB1" &
    x"860E5E0A_5A3E2AB3_771FE71C_4E3D06FA_2965DCB9_99E71D0F" &
    x"803E89D6_5266C825_2E4CC978_9C10B36A_C6150EBA_94E2EA78" &
    x"A5FC3C53_1E0A2DF4_F2F74EA7_361D2B3D_1939260F_19C27960" &
    x"5223A708_F71312B6_EBADFE6E_EAC31F66_E3BC4595_A67BC883" &
    x"B17F37D1_018CFF28_C332DDEF_BE6C5AA5_65582185_68AB9802" &
    x"EECEA50F_DB2F953B_2AEF7DAD_5B6E2F84_1521B628_29076170" &
    x"ECDD4775_619F1510_13CCA830_EB61BD96_0334FE1E_AA0363CF" &
    x"B5735C90_4C70A239_D59E9E0B_CBAADE14_EECC86BC_60622CA7" &
    x"9CAB5CAB_B2F3846E_648B1EAF_19BDF0CA_A02369B9_655ABB50" &
    x"40685A32_3C2AB4B3_319EE9D5_C021B8F7_9B540B19_875FA099" &
    x"95F7997E_623D7DA8_F837889A_97E32D77_11ED935F_16681281" &
    x"0E358829_C7E61FD6_96DEDFA1_7858BA99_57F584A5_1B227263" &
    x"9B83C3FF_1AC24696_CDB30AEB_532E3054_8FD948E4_6DBC3128" &
    x"58EBF2EF_34C6FFEA_FE28ED61_EE7C3C73_5D4A14D9_E864B7E3" &
    x"42105D14_203E13E0_45EEE2B6_A3AAABEA_DB6C4F15_FACB4FD0" &
    x"C742F442_EF6ABBB5_654F3B1D_41CD2105_D81E799E_86854DC7" &
    x"E44B476A_3D816250_CF62A1F2_5B8D2646_FC8883A0_C1C7B6A3" &
    x"7F1524C3_69CB7492_47848A0B_5692B285_095BBF00_AD19489D" &
    x"1462B174_23820E00_58428D2A_0C55F5EA_1DADF43E_233F7061" &
    x"3372F092_8D937E41_D65FECF1_6C223BDB_7CDE3759_CBEE7460" &
    x"4085F2A7_CE77326E_A6078084_19F8509E_E8EFD855_61D99735" &
    x"A969A7AA_C50C06C2_5A04ABFC_800BCADC_9E447A2E_C3453484" &
    x"FDD56705_0E1E9EC9_DB73DBD3_105588CD_675FDA79_E3674340" &
    x"C5C43465_713E38D8_3D28F89E_F16DFF20_153E21E7_8FB03D4A" &
    x"E6E39F2B_DB83ADF7";
    
    constant SBOX23_INIT_VEC : std_logic_vector(16383 downto 0) :=
    x"E93D5A68_948140F7_F64C261C_94692934_411520F7_7602D4F7" &
    x"BCF46B2E_D4A20068_D4082471_3320F46A_43B7D4B7_500061AF" &
    x"1E39F62E_97244546_14214F74_BF8B8840_4D95FC1D_96B591AF" &
    x"70F4DDD3_66A02F45_BFBC09EC_03BD9785_7FAC6DD0_31CB8504" &
    x"96EB27B3_55FD3941_DA2547E6_ABCA0A9A_28507825_530429F4" &
    x"0A2C86DA_E9B66DFB_68DC1462_D7486900_680EC0A4_27A18DEE" &
    x"4F3FFEA2_E887AD8C_B58CE006_7AF4D6B6_AACE1E7C_D3375FEC" &
    x"CE78A399_406B2A42_20FE9E35_D9F385B9_EE39D7AB_3B124E8B" &
    x"1DC9FAF7_4B6D1856_26A36631_EAE397B2_3A6EFA74_DD5B4332" &
    x"6841E7F7_CA7820FB_FB0AF54E_D8FEB397_454056AC_BA489527" &
    x"55533A3A_20838D87_FE6BA9B7_D096954B_55A867BC_A1159A58" &
    x"CCA92963_99E1DB33_A62A4A56_3F3125F9_5EF47E1C_9029317C" &
    x"FDF8E802_04272F70_80BB155C_05282CE3_95C11548_E4C66D22" &
    x"48C1133F_C70F86DC_07F9C9EE_41041F0F_404779A4_5D886E17" &
    x"325F51EB_D59BC0D1_F2BCC18F_41113564_257B7834_602A9C60" &
    x"DFF8E8A3_1F636C1B_0E12B4C2_02E1329E_AF664FD1_CAD18115" &
    x"6B2395E0_333E92E1_3B240B62_EEBEB922_85B2A20E_E6BA0D99" &
    x"DE720C8C_2DA2F728_D0127845_95B794FD_647D0862_E7CCF5F0" &
    x"5449A36F_877D48FA_C39DFD27_F33E8D1E_0A476341_992EFF74" &
    x"3A6F6EAB_F4F8FD37_A812DC60_A1EBDDF8_991BE14C_DB6E6B0D" &
    x"C67B5510_6D672C37_2765D43B_DCD0E804_F1290DC7_CC00FFA3" &
    x"B5390F92_690FED0B_667B9FFB_CEDB7D9C_A091CF0B_D9155EA3" &
    x"BB132F88_515BAD24_7B9479BF_763BD6EB_37392EB3_CC115979" &
    x"8026E297_F42E312D_6842ADA7_C66A2B3B_12754CCC_782EF11C" &
    x"6A124237_B79251E7_06A1BBE6_4BFB6350_1A6B1018_11CAEDFA" &
    x"3D25BDD8_E2E1C3C9_44421659_0A121386_D90CEC6E_D5ABEA2A" &
    x"64AF674E_DA86A85F_BEBFE988_64E4C3FE_9DBC8057_F0F7C086" &
    x"60787BF8_6003604D_D1FD8346_F6381FB0_7745AE04_D736FCCC" &
    x"83426B33_F01EAB71_B0804187_3C005E5F_77A057BE_BDE8AE24" &
    x"55464299_BF582E61_4E58F48F_F2DDFDA2_F474EF38_8789BDC2" &
    x"5366F9C3_C8B38E74_B475F255_46FCD9B9_7AEB2661_8B1DDF84" &
    x"846A0E79_915F95E2_466E598E_20B45770_8CD55591_C902DE4C" &
    x"B90BACE1_BB8205D0_11A86248_7574A99E_B77F19B6_E0A9DC09" &
    x"662D09A1_C4324633_E85A1F02_09F0BE8C_4A99A025_1D6EFE10" &
    x"1AB93D1D_0BA5A4DF_A186F20F_2868F169_DCB7DA83_573906FE" &
    x"A1E2CE9B_4FCD7F52_50115E01_A70683FA_A002B5C4_0DE6D027" &
    x"9AF88C27_773F8641_C3604C06_61A806B5_F0177A28_C0F586E0" &
    x"006058AA_30DC7D62_11E69ED7_2338EA63_53C2DD94_C2C21634" &
    x"BBCBEE56_90BCB6DE_EBFC7DA1_CE591D76_6F05E409_4B7C0188" &
    x"39720A3D_7C927C24_86E3725F_724D9DB9_1AC15BB4_D39EB8FC" &
    x"ED545578_08FCA5B5_D83D7CD3_4DAD0FC4_1E50EF5E_B161E6F8" &
    x"A28514D9_6C51133C_6FD5C7E7_56E14EC4_362ABFCE_DDC6C837" &
    x"D79A3234_92638212_670EFA8E_406000E0_3A39CE37_D3FAF5CF" &
    x"ABC27737_5AC52D1B_5CB0679E_4FA33742_D3822740_99BC9BBE" &
    x"D5118E9D_BF0F7315_D62D1C7E_C700C47B_B78C1B6B_21A19045" &
    x"B26EB1BE_6A366EB4_5748AB2F_BC946E79_C6A376D2_6549C2C8" &
    x"530FF8EE_468DDE7D_D5730A1D_4CD04DC6_2939BBDB_A9BA4650" &
    x"AC9526E8_BE5EE304_A1FAD5F0_6A2D519A_63EF8CE2_9A86EE22" &
    x"C089C2B8_43242EF6_A51E03AA_9CF2D0A4_83C061BA_9BE96A4D" &
    x"8FE51550_BA645BD6_2826A2F9_A73A3AE1_4BA99586_EF5562E9" &
    x"C72FEFD3_F752F7DA_3F046F69_77FA0A59_80E4A915_87B08601" &
    x"9B09E6AD_3B3EE593_E990FD5A_9E34D797_2CF0B7D9_022B8B51" &
    x"96D5AC3A_017DA67D_D1CF3ED6_7C7D2D28_1F9F25CF_ADF2B89B" &
    x"5AD6B472_5A88F54C_E029AC71_E019A5E6_47B0ACFD_ED93FA9B" &
    x"E8D3C48D_283B57CC_F8D56629_79132E28_785F0191_ED756055" &
    x"F7960E44_E3D35E8C_15056DD4_88F46DBA_03A16125_0564F0BD" &
    x"C3EB9E15_3C9057A2_97271AEC_A93A072A_1B3F6D9B_1E6321F5" &
    x"F59C66FB_26DCF319_7533D928_B155FDF5_03563482_8ABA3CBB" &
    x"28517711_C20AD9F8_ABCC5167_CCAD925F_4DE81751_3830DC8E" &
    x"379D5862_9320F991_EA7A90C2_FB3E7BCE_5121CE64_774FBE32" &
    x"A8B6E37E_C3293D46_48DE5369_6413E680_A2AE0810_DD6DB224" &
    x"69852DFD_09072166_B39A460A_6445C0DD_586CDECF_1C20C8AE" &
    x"5BBEF7DD_1B588D40_CCD2017F_6BB4E3BB_DDA26A7E_3A59FF45" &
    x"3E350A44_BCB4CDD5_72EACEA8_FA6484BB_8D6612AE_BF3C6F47" &
    x"D29BE463_542F5D9E_AEC2771B_F64E6370_740E0D8D_E75B1357" &
    x"F8721671_AF537D5D_4040CB08_4EB4E2CC_34D2466A_0115AF84" &
    x"E1B00428_95983A1D_06B89FB4_CE6EA048_6F3F3B82_3520AB82" &
    x"011A1D4B_277227F8_611560B1_E7933FDC_BB3A792B_344525BD" &
    x"A08839E1_51CE794B_2F32C9B7_A01FBAC9_E01CC87E_BCC7D1F6" &
    x"CF0111C3_A1E8AAC7_1A908749_D44FBD9A_D0DADECB_D50ADA38" &
    x"0339C32A_C6913667_8DF9317C_E0B12B4F_F79E59B7_43F5BB3A" &
    x"F2D519FF_27D9459C_BF97222C_15E6FC2A_0F91FC71_9B941525" &
    x"FAE59361_CEB69CEB_C2A86459_12BAA8D1_B6C1075E_E3056A0C" &
    x"10D25065_CB03A442_E0EC6E0E_1698DB3B_4C98A0BE_3278E964" &
    x"9F1F9532_E0D392DF_D3A0342B_8971F21E_1B0A7441_4BA3348C" &
    x"C5BE7120_C37632D8_DF359F8D_9B992F2E_E60B6F47_0FE3F11D" &
    x"E54CDA54_1EDAD891_CE6279CF_CD3E7E6F_1618B166_FD2C1D05" &
    x"848FD2C5_F6FB2299_F523F357_A6327623_93A83531_56CCCD02" &
    x"ACF08162_5A75EBB5_6E163697_88D273CC_DE966292_81B949D0" &
    x"4C50901B_71C65614_E6C6C7BD_327A140A_45E1D006_C3F27B9A" &
    x"C9AA53FD_62A80F00_BB25BFE2_35BDD2F6_71126905_B2040222" &
    x"B6CBCF7C_CD769C2B_53113EC0_1640E3D3_38ABBD60_2547ADF0" &
    x"BA38209C_F746CE76_77AFA1C5_20756060_85CBFE4E_8AE88DD8" &
    x"7AAAF9B0_4CF9AA7E_1948C25C_02FB8A8C_01C36AE4_D6EBE1F9" &
    x"90D4F869_A65CDEA0_3F09252D_C208E69F_B74E6132_CE77E25B" &
    x"578FDFE3_3AC372E6";
end package pkg_sbox_init;